module double_threshold_unit (); 



endmodule 


