module peripheral (
    input wire clk,
    input wire reset_n
); endmodule 



//Module to output the output of the Image Detector

