module hysterisis_unit (

); 






endmodule 


